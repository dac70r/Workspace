
module my_timer (
	clk_clk,
	led_export);	

	input		clk_clk;
	output		led_export;
endmodule
