
module PLL_complete (
	clk_clk,
	reset_reset_n,
	to_outside_led);	

	input		clk_clk;
	input		reset_reset_n;
	output		to_outside_led;
endmodule
