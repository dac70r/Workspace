
module My_First_NIOS_II_Platform_Designer (
	clk_clk,
	gpio_external_connection_export);	

	input		clk_clk;
	output	[7:0]	gpio_external_connection_export;
endmodule
