
/* Top level HDL module that instatiates the 
	embedded system
*/

module component_tutorial (CLOCK_50, KEY, HEX0, HEX1, HEX2, HEX3);

input CLOCK_50;
input [0:0] KEY;
output [0:6] HEX0, HEX1, HEX2, HEX3;

wire [15:0] to_HEX;

unsaved_unfinished U0 (
.clk_clk(CLOCK_50), .resetn_reset_n(KEY[0]), .to_hex_export(to_HEX) );

hex7seg h0(to_HEX[3:0], HEX0);
hex7seg h1(to_HEX[7:4], HEX1);
hex7seg h2(to_HEX[11:8], HEX2);
hex7seg h3(to_HEX[15:12], HEX3);

endmodule