
module My_First_NIOS_II_Platform_Designer (
	clk_clk,
	gpio_external_connection_export,
	reset_reset_n);	

	input		clk_clk;
	output	[7:0]	gpio_external_connection_export;
	input		reset_reset_n;
endmodule
