// My_First_NIOS_II_Platform_Designer.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module My_First_NIOS_II_Platform_Designer (
		input  wire       clk_clk,                         //                      clk.clk
		output wire [7:0] gpio_external_connection_export  // gpio_external_connection.export
	);

	wire         hellonios_debug_reset_request_reset;                     // HelloNios:debug_reset_request -> rst_controller:reset_in0
	wire  [31:0] hellonios_data_master_readdata;                          // mm_interconnect_0:HelloNios_data_master_readdata -> HelloNios:d_readdata
	wire         hellonios_data_master_waitrequest;                       // mm_interconnect_0:HelloNios_data_master_waitrequest -> HelloNios:d_waitrequest
	wire         hellonios_data_master_debugaccess;                       // HelloNios:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:HelloNios_data_master_debugaccess
	wire  [13:0] hellonios_data_master_address;                           // HelloNios:d_address -> mm_interconnect_0:HelloNios_data_master_address
	wire   [3:0] hellonios_data_master_byteenable;                        // HelloNios:d_byteenable -> mm_interconnect_0:HelloNios_data_master_byteenable
	wire         hellonios_data_master_read;                              // HelloNios:d_read -> mm_interconnect_0:HelloNios_data_master_read
	wire         hellonios_data_master_write;                             // HelloNios:d_write -> mm_interconnect_0:HelloNios_data_master_write
	wire  [31:0] hellonios_data_master_writedata;                         // HelloNios:d_writedata -> mm_interconnect_0:HelloNios_data_master_writedata
	wire  [31:0] hellonios_instruction_master_readdata;                   // mm_interconnect_0:HelloNios_instruction_master_readdata -> HelloNios:i_readdata
	wire         hellonios_instruction_master_waitrequest;                // mm_interconnect_0:HelloNios_instruction_master_waitrequest -> HelloNios:i_waitrequest
	wire  [13:0] hellonios_instruction_master_address;                    // HelloNios:i_address -> mm_interconnect_0:HelloNios_instruction_master_address
	wire         hellonios_instruction_master_read;                       // HelloNios:i_read -> mm_interconnect_0:HelloNios_instruction_master_read
	wire         mm_interconnect_0_debug_avalon_jtag_slave_chipselect;    // mm_interconnect_0:DEBUG_avalon_jtag_slave_chipselect -> DEBUG:av_chipselect
	wire  [31:0] mm_interconnect_0_debug_avalon_jtag_slave_readdata;      // DEBUG:av_readdata -> mm_interconnect_0:DEBUG_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_debug_avalon_jtag_slave_waitrequest;   // DEBUG:av_waitrequest -> mm_interconnect_0:DEBUG_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_debug_avalon_jtag_slave_address;       // mm_interconnect_0:DEBUG_avalon_jtag_slave_address -> DEBUG:av_address
	wire         mm_interconnect_0_debug_avalon_jtag_slave_read;          // mm_interconnect_0:DEBUG_avalon_jtag_slave_read -> DEBUG:av_read_n
	wire         mm_interconnect_0_debug_avalon_jtag_slave_write;         // mm_interconnect_0:DEBUG_avalon_jtag_slave_write -> DEBUG:av_write_n
	wire  [31:0] mm_interconnect_0_debug_avalon_jtag_slave_writedata;     // mm_interconnect_0:DEBUG_avalon_jtag_slave_writedata -> DEBUG:av_writedata
	wire  [31:0] mm_interconnect_0_hellonios_debug_mem_slave_readdata;    // HelloNios:debug_mem_slave_readdata -> mm_interconnect_0:HelloNios_debug_mem_slave_readdata
	wire         mm_interconnect_0_hellonios_debug_mem_slave_waitrequest; // HelloNios:debug_mem_slave_waitrequest -> mm_interconnect_0:HelloNios_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_hellonios_debug_mem_slave_debugaccess; // mm_interconnect_0:HelloNios_debug_mem_slave_debugaccess -> HelloNios:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_hellonios_debug_mem_slave_address;     // mm_interconnect_0:HelloNios_debug_mem_slave_address -> HelloNios:debug_mem_slave_address
	wire         mm_interconnect_0_hellonios_debug_mem_slave_read;        // mm_interconnect_0:HelloNios_debug_mem_slave_read -> HelloNios:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_hellonios_debug_mem_slave_byteenable;  // mm_interconnect_0:HelloNios_debug_mem_slave_byteenable -> HelloNios:debug_mem_slave_byteenable
	wire         mm_interconnect_0_hellonios_debug_mem_slave_write;       // mm_interconnect_0:HelloNios_debug_mem_slave_write -> HelloNios:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_hellonios_debug_mem_slave_writedata;   // mm_interconnect_0:HelloNios_debug_mem_slave_writedata -> HelloNios:debug_mem_slave_writedata
	wire         mm_interconnect_0_sram_s1_chipselect;                    // mm_interconnect_0:SRAM_s1_chipselect -> SRAM:chipselect
	wire  [31:0] mm_interconnect_0_sram_s1_readdata;                      // SRAM:readdata -> mm_interconnect_0:SRAM_s1_readdata
	wire   [9:0] mm_interconnect_0_sram_s1_address;                       // mm_interconnect_0:SRAM_s1_address -> SRAM:address
	wire   [3:0] mm_interconnect_0_sram_s1_byteenable;                    // mm_interconnect_0:SRAM_s1_byteenable -> SRAM:byteenable
	wire         mm_interconnect_0_sram_s1_write;                         // mm_interconnect_0:SRAM_s1_write -> SRAM:write
	wire  [31:0] mm_interconnect_0_sram_s1_writedata;                     // mm_interconnect_0:SRAM_s1_writedata -> SRAM:writedata
	wire         mm_interconnect_0_sram_s1_clken;                         // mm_interconnect_0:SRAM_s1_clken -> SRAM:clken
	wire         mm_interconnect_0_gpio_s1_chipselect;                    // mm_interconnect_0:GPIO_s1_chipselect -> GPIO:chipselect
	wire  [31:0] mm_interconnect_0_gpio_s1_readdata;                      // GPIO:readdata -> mm_interconnect_0:GPIO_s1_readdata
	wire   [1:0] mm_interconnect_0_gpio_s1_address;                       // mm_interconnect_0:GPIO_s1_address -> GPIO:address
	wire         mm_interconnect_0_gpio_s1_write;                         // mm_interconnect_0:GPIO_s1_write -> GPIO:write_n
	wire  [31:0] mm_interconnect_0_gpio_s1_writedata;                     // mm_interconnect_0:GPIO_s1_writedata -> GPIO:writedata
	wire         mm_interconnect_0_timer_s1_chipselect;                   // mm_interconnect_0:TIMER_s1_chipselect -> TIMER:chipselect
	wire  [15:0] mm_interconnect_0_timer_s1_readdata;                     // TIMER:readdata -> mm_interconnect_0:TIMER_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_s1_address;                      // mm_interconnect_0:TIMER_s1_address -> TIMER:address
	wire         mm_interconnect_0_timer_s1_write;                        // mm_interconnect_0:TIMER_s1_write -> TIMER:write_n
	wire  [15:0] mm_interconnect_0_timer_s1_writedata;                    // mm_interconnect_0:TIMER_s1_writedata -> TIMER:writedata
	wire         irq_mapper_receiver0_irq;                                // DEBUG:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                // TIMER:irq -> irq_mapper:receiver1_irq
	wire  [31:0] hellonios_irq_irq;                                       // irq_mapper:sender_irq -> HelloNios:irq
	wire         rst_controller_reset_out_reset;                          // rst_controller:reset_out -> [DEBUG:rst_n, GPIO:reset_n, HelloNios:reset_n, SRAM:reset, TIMER:reset_n, irq_mapper:reset, mm_interconnect_0:HelloNios_reset_reset_bridge_in_reset_reset, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                      // rst_controller:reset_req -> [HelloNios:reset_req, SRAM:reset_req, rst_translator:reset_req_in]

	My_First_NIOS_II_Platform_Designer_DEBUG debug (
		.clk            (clk_clk),                                               //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_debug_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_debug_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_debug_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_debug_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_debug_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_debug_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_debug_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                               //               irq.irq
	);

	My_First_NIOS_II_Platform_Designer_GPIO gpio (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_gpio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_gpio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_gpio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_gpio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_gpio_s1_readdata),   //                    .readdata
		.out_port   (gpio_external_connection_export)       // external_connection.export
	);

	My_First_NIOS_II_Platform_Designer_HelloNios hellonios (
		.clk                                 (clk_clk),                                                 //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                         //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                      //                          .reset_req
		.d_address                           (hellonios_data_master_address),                           //               data_master.address
		.d_byteenable                        (hellonios_data_master_byteenable),                        //                          .byteenable
		.d_read                              (hellonios_data_master_read),                              //                          .read
		.d_readdata                          (hellonios_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (hellonios_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (hellonios_data_master_write),                             //                          .write
		.d_writedata                         (hellonios_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (hellonios_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (hellonios_instruction_master_address),                    //        instruction_master.address
		.i_read                              (hellonios_instruction_master_read),                       //                          .read
		.i_readdata                          (hellonios_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (hellonios_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (hellonios_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (hellonios_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_hellonios_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_hellonios_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_hellonios_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_hellonios_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_hellonios_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_hellonios_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_hellonios_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_hellonios_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                         // custom_instruction_master.readra
	);

	My_First_NIOS_II_Platform_Designer_SRAM sram (
		.clk        (clk_clk),                              //   clk1.clk
		.address    (mm_interconnect_0_sram_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_sram_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_sram_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_sram_s1_write),      //       .write
		.readdata   (mm_interconnect_0_sram_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_sram_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_sram_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),       // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),   //       .reset_req
		.freeze     (1'b0)                                  // (terminated)
	);

	My_First_NIOS_II_Platform_Designer_TIMER timer (
		.clk        (clk_clk),                               //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       // reset.reset_n
		.address    (mm_interconnect_0_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)               //   irq.irq
	);

	My_First_NIOS_II_Platform_Designer_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                               (clk_clk),                                                 //                             clk_0_clk.clk
		.HelloNios_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                          // HelloNios_reset_reset_bridge_in_reset.reset
		.HelloNios_data_master_address               (hellonios_data_master_address),                           //                 HelloNios_data_master.address
		.HelloNios_data_master_waitrequest           (hellonios_data_master_waitrequest),                       //                                      .waitrequest
		.HelloNios_data_master_byteenable            (hellonios_data_master_byteenable),                        //                                      .byteenable
		.HelloNios_data_master_read                  (hellonios_data_master_read),                              //                                      .read
		.HelloNios_data_master_readdata              (hellonios_data_master_readdata),                          //                                      .readdata
		.HelloNios_data_master_write                 (hellonios_data_master_write),                             //                                      .write
		.HelloNios_data_master_writedata             (hellonios_data_master_writedata),                         //                                      .writedata
		.HelloNios_data_master_debugaccess           (hellonios_data_master_debugaccess),                       //                                      .debugaccess
		.HelloNios_instruction_master_address        (hellonios_instruction_master_address),                    //          HelloNios_instruction_master.address
		.HelloNios_instruction_master_waitrequest    (hellonios_instruction_master_waitrequest),                //                                      .waitrequest
		.HelloNios_instruction_master_read           (hellonios_instruction_master_read),                       //                                      .read
		.HelloNios_instruction_master_readdata       (hellonios_instruction_master_readdata),                   //                                      .readdata
		.DEBUG_avalon_jtag_slave_address             (mm_interconnect_0_debug_avalon_jtag_slave_address),       //               DEBUG_avalon_jtag_slave.address
		.DEBUG_avalon_jtag_slave_write               (mm_interconnect_0_debug_avalon_jtag_slave_write),         //                                      .write
		.DEBUG_avalon_jtag_slave_read                (mm_interconnect_0_debug_avalon_jtag_slave_read),          //                                      .read
		.DEBUG_avalon_jtag_slave_readdata            (mm_interconnect_0_debug_avalon_jtag_slave_readdata),      //                                      .readdata
		.DEBUG_avalon_jtag_slave_writedata           (mm_interconnect_0_debug_avalon_jtag_slave_writedata),     //                                      .writedata
		.DEBUG_avalon_jtag_slave_waitrequest         (mm_interconnect_0_debug_avalon_jtag_slave_waitrequest),   //                                      .waitrequest
		.DEBUG_avalon_jtag_slave_chipselect          (mm_interconnect_0_debug_avalon_jtag_slave_chipselect),    //                                      .chipselect
		.GPIO_s1_address                             (mm_interconnect_0_gpio_s1_address),                       //                               GPIO_s1.address
		.GPIO_s1_write                               (mm_interconnect_0_gpio_s1_write),                         //                                      .write
		.GPIO_s1_readdata                            (mm_interconnect_0_gpio_s1_readdata),                      //                                      .readdata
		.GPIO_s1_writedata                           (mm_interconnect_0_gpio_s1_writedata),                     //                                      .writedata
		.GPIO_s1_chipselect                          (mm_interconnect_0_gpio_s1_chipselect),                    //                                      .chipselect
		.HelloNios_debug_mem_slave_address           (mm_interconnect_0_hellonios_debug_mem_slave_address),     //             HelloNios_debug_mem_slave.address
		.HelloNios_debug_mem_slave_write             (mm_interconnect_0_hellonios_debug_mem_slave_write),       //                                      .write
		.HelloNios_debug_mem_slave_read              (mm_interconnect_0_hellonios_debug_mem_slave_read),        //                                      .read
		.HelloNios_debug_mem_slave_readdata          (mm_interconnect_0_hellonios_debug_mem_slave_readdata),    //                                      .readdata
		.HelloNios_debug_mem_slave_writedata         (mm_interconnect_0_hellonios_debug_mem_slave_writedata),   //                                      .writedata
		.HelloNios_debug_mem_slave_byteenable        (mm_interconnect_0_hellonios_debug_mem_slave_byteenable),  //                                      .byteenable
		.HelloNios_debug_mem_slave_waitrequest       (mm_interconnect_0_hellonios_debug_mem_slave_waitrequest), //                                      .waitrequest
		.HelloNios_debug_mem_slave_debugaccess       (mm_interconnect_0_hellonios_debug_mem_slave_debugaccess), //                                      .debugaccess
		.SRAM_s1_address                             (mm_interconnect_0_sram_s1_address),                       //                               SRAM_s1.address
		.SRAM_s1_write                               (mm_interconnect_0_sram_s1_write),                         //                                      .write
		.SRAM_s1_readdata                            (mm_interconnect_0_sram_s1_readdata),                      //                                      .readdata
		.SRAM_s1_writedata                           (mm_interconnect_0_sram_s1_writedata),                     //                                      .writedata
		.SRAM_s1_byteenable                          (mm_interconnect_0_sram_s1_byteenable),                    //                                      .byteenable
		.SRAM_s1_chipselect                          (mm_interconnect_0_sram_s1_chipselect),                    //                                      .chipselect
		.SRAM_s1_clken                               (mm_interconnect_0_sram_s1_clken),                         //                                      .clken
		.TIMER_s1_address                            (mm_interconnect_0_timer_s1_address),                      //                              TIMER_s1.address
		.TIMER_s1_write                              (mm_interconnect_0_timer_s1_write),                        //                                      .write
		.TIMER_s1_readdata                           (mm_interconnect_0_timer_s1_readdata),                     //                                      .readdata
		.TIMER_s1_writedata                          (mm_interconnect_0_timer_s1_writedata),                    //                                      .writedata
		.TIMER_s1_chipselect                         (mm_interconnect_0_timer_s1_chipselect)                    //                                      .chipselect
	);

	My_First_NIOS_II_Platform_Designer_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.sender_irq    (hellonios_irq_irq)               //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (hellonios_debug_reset_request_reset), // reset_in0.reset
		.clk            (clk_clk),                             //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),      // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),  //          .reset_req
		.reset_req_in0  (1'b0),                                // (terminated)
		.reset_in1      (1'b0),                                // (terminated)
		.reset_req_in1  (1'b0),                                // (terminated)
		.reset_in2      (1'b0),                                // (terminated)
		.reset_req_in2  (1'b0),                                // (terminated)
		.reset_in3      (1'b0),                                // (terminated)
		.reset_req_in3  (1'b0),                                // (terminated)
		.reset_in4      (1'b0),                                // (terminated)
		.reset_req_in4  (1'b0),                                // (terminated)
		.reset_in5      (1'b0),                                // (terminated)
		.reset_req_in5  (1'b0),                                // (terminated)
		.reset_in6      (1'b0),                                // (terminated)
		.reset_req_in6  (1'b0),                                // (terminated)
		.reset_in7      (1'b0),                                // (terminated)
		.reset_req_in7  (1'b0),                                // (terminated)
		.reset_in8      (1'b0),                                // (terminated)
		.reset_req_in8  (1'b0),                                // (terminated)
		.reset_in9      (1'b0),                                // (terminated)
		.reset_req_in9  (1'b0),                                // (terminated)
		.reset_in10     (1'b0),                                // (terminated)
		.reset_req_in10 (1'b0),                                // (terminated)
		.reset_in11     (1'b0),                                // (terminated)
		.reset_req_in11 (1'b0),                                // (terminated)
		.reset_in12     (1'b0),                                // (terminated)
		.reset_req_in12 (1'b0),                                // (terminated)
		.reset_in13     (1'b0),                                // (terminated)
		.reset_req_in13 (1'b0),                                // (terminated)
		.reset_in14     (1'b0),                                // (terminated)
		.reset_req_in14 (1'b0),                                // (terminated)
		.reset_in15     (1'b0),                                // (terminated)
		.reset_req_in15 (1'b0)                                 // (terminated)
	);

endmodule
