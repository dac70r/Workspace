
module EtherCAT (
	clk_clk,
	led_export,
	reset_reset_n,
	timer_export);	

	input		clk_clk;
	output		led_export;
	input		reset_reset_n;
	output		timer_export;
endmodule
